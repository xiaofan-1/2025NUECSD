`timescale 1ns / 1ps

module arp_ctrl(
    input   wire            clk             ,
    input   wire            rst_n           ,
    input   wire            key             ,
    input   wire            arp_rx_op       ,
    input   wire            arp_rx_done     ,
    output  reg             arp_tx_en       ,
    output  reg             arp_tx_op        //1:�����/0:Ӧ���
    );
    
always @(posedge clk) begin
    if(!rst_n) begin
        arp_tx_en <= 0;
        arp_tx_op <= 0;
    end
    else if(key) begin //���������
        arp_tx_en <= 1;
        arp_tx_op <= 1;
    end
    else if(arp_rx_op == 1 && arp_rx_done) begin //���յ������������Ӧ���
        arp_tx_en <= 1;
        arp_tx_op <= 0;
    end
    else if(arp_rx_op == 0 && arp_rx_done) begin //���յ�Ӧ�����������
        arp_tx_en <= 0;
        arp_tx_op <= 0;
    end
    else begin
        arp_tx_en <= 0;
        arp_tx_op <= arp_tx_op;
    end
end
endmodule
