`timescale 1ns / 1ps

module image_data #(
    parameter	H_PIXEL = 16'd1280,//�ֱ���Ϊ1280*720
    parameter	V_PIXEL = 16'd720  //һ��udp������1280�ֽڣ���Ҫ����1440��
)(
    input   wire            clk                 ,
    input   wire            rst_n               ,
    
    input   wire    [7:0]   cam_data            ,//ddr����ͷ����
    input   wire            udp_data_start      ,//��ʼִ�б�ģ���ź�
    input   wire            udp_tx_done         ,//��̫��������һ���������ź�
    input   wire            rf_rd_req           ,//ddr��fifo��Ϊ���ź�
    input   wire            udp_data_valid      ,//udp������Ч�ź�
   
    output  wire            rf_rd_en            ,//ddr��fifoʹ��
    output  reg     [7:0]   image_data          ,//��װ�õ�ͼ������
    output  reg             udp_tx_data_start   ,//��̫����ʼ�����ź�
    output  reg     [15:0]  image_data_num       //��̫���������ݸ���
    );
	
localparam
    CNT_PACKET_WAIT = 28'd10,
    CNT_FRAME_WAIT = 28'd10;
    
localparam
    HEAD     =   32'h53_5a_48_59 ,//��ͷ
    ADDR     =   8'h00           ,//�豸��ַ
    CMD      =   8'h02           ,//ָ��
    CRC      =   16'h7C_0B       ;//CRC-16У�飺�ر���λ��У�飬����д����ֵ

localparam
    IDLE        = 6'b000_001,                               
    HEAD_PACKET = 6'b000_010,//��һ�����ݣ�������ͷ    
	DATA_STARTE = 6'b100_001,
    DATA_PACKET = 6'b000_100,//ͼ������
	LAST_STARTE = 6'b100_010,
    LAST_PACKET = 6'b001_000,//���һ������
    PACKET_WAIT = 6'b010_000,//���������꣬�ȴ�ʱ��
    FRAME_WAIT  = 6'b100_000;//һ֡���ݷ����꣬�ȴ�ʱ��

reg     [5:0]   curr_state;
reg     [5:0]   next_state;
reg     [27:0]  cnt_packet;//�����ȴ�ʱ�����
reg     [27:0]  cnt_frame;//��֡�ȴ�ʱ�����
//reg     [10:0]  cnt_v;//
reg     [10:0]  cnt_h;//һ֡ͼ����udp���ĸ���
reg     [10:0]  cnt_data;//�������ݸ���������2�ֽ�

reg             udp_data_start_reg;
reg             udp_data_valid_reg;

localparam TOTAL_BYTES_VALUE = H_PIXEL*V_PIXEL*2 + 4 + 1 + 4 + 1 + 2;//��������ʾ�Ӱ�ͷ��У����������ݳ��ȣ���λΪ�ֽ�   00_1c_20_0c   00_09_60_0c
                         //(1280*720*2)(ͼ������) + 4(��ͷ) + 1(�豸��ַ) + 4(������) + 1(ָ���ֽ�) + 2(У���ֽ�)

// ����һ�� wire����ʹ��ƴ�Ӳ����������ֽڷ�ת���õ�С����
wire	[31:0]	DATA_NUM ;
assign DATA_NUM = {TOTAL_BYTES_VALUE[7:0],   // Byte 0 (LSB)
                   TOTAL_BYTES_VALUE[15:8],  // Byte 1
                   TOTAL_BYTES_VALUE[23:16], // Byte 2
                   TOTAL_BYTES_VALUE[31:24]};// Byte 3 (MSB)
				   
wire	[15:0]	h_num;
wire	[15:0]	v_num;
assign	h_num = (H_PIXEL <= 16'd736) ? H_PIXEL*2 : H_PIXEL;
assign	v_num = (H_PIXEL <= 16'd736) ? V_PIXEL : V_PIXEL*2;

//----------------------------state_one----------------------
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        curr_state <= IDLE;
    else
        curr_state <= next_state;
end

//----------------------------state_two----------------------
always @(*) begin
    if(!rst_n)
        next_state = IDLE;
    else begin
        case(curr_state)
            IDLE       :begin
                if(rf_rd_req && udp_data_start)
                    next_state = HEAD_PACKET;
                else
                    next_state = curr_state;
            end
            HEAD_PACKET:begin//��һ�����ݣ�������ͷ
                if(udp_tx_done)
                    next_state = PACKET_WAIT;
                else
                    next_state = curr_state;
            end
			DATA_STARTE:begin
                if(rf_rd_req && udp_data_start)
                    next_state = DATA_PACKET;
                else
                    next_state = curr_state;
            end
            DATA_PACKET:begin//ͼ������
                if(udp_tx_done)
                    next_state = PACKET_WAIT;
                else
                    next_state = curr_state;
            end
			LAST_STARTE:begin
                if(rf_rd_req && udp_data_start)
                    next_state = LAST_PACKET;
                else
                    next_state = curr_state;
            end
            LAST_PACKET: begin//���һ������
                if(udp_tx_done)
                    next_state = IDLE;
                else
                    next_state = curr_state;
            end
            PACKET_WAIT: begin//���������꣬�ȴ�ʱ��
                if(cnt_h < v_num - 16'd1)
                    next_state = DATA_STARTE;
                else if(cnt_h == v_num - 16'd1)
                    next_state = LAST_STARTE;
                else
                    next_state = curr_state;
            end
            FRAME_WAIT : begin//һ֡���ݷ����꣬�ȴ�ʱ��
                if(cnt_frame == CNT_FRAME_WAIT)
                    next_state = IDLE;
                else
                    next_state = curr_state;
            end
            default:next_state = IDLE;
        endcase
    end
end
//-----------------------------��ʼִ�б�ģ���ź�------------------------
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        udp_data_start_reg <= 1'b0;
    else if(udp_data_start)
        udp_data_start_reg <= 1'b1;
    else
        udp_data_start_reg <= udp_data_start_reg;
end
//----------------------------����udp_data_valid----------------------
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        udp_data_valid_reg <= 1'b0;
    else
        udp_data_valid_reg <= udp_data_valid;
end
//----------------------------�������ݵȴ�ʱ��----------------------
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        cnt_packet <= 28'd0;
    else if((curr_state == IDLE || curr_state == PACKET_WAIT) && udp_data_start_reg) begin
        if(cnt_packet == CNT_PACKET_WAIT)
            cnt_packet <= 28'd0;
        else
            cnt_packet <= cnt_packet + 28'd1;
    end
    else
        cnt_packet <= 28'd0;
end
//----------------------------��֡���ݵȴ�ʱ��----------------------
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        cnt_frame <= 28'd0;
    else if(curr_state == FRAME_WAIT) begin
        if(cnt_frame == CNT_FRAME_WAIT)
            cnt_frame <= 28'd0;
        else
            cnt_frame <= cnt_frame + 1;
    end
    else
        cnt_frame <= 28'd0;
end
//----------------------------�������ݼ���----------------------
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        cnt_data <= 11'd0;
    else if(curr_state == HEAD_PACKET || curr_state == DATA_PACKET || curr_state == LAST_PACKET) begin
        if(udp_data_valid_reg)
            cnt_data <= cnt_data + 1;
        else
            cnt_data <= cnt_data;
    end
    else
        cnt_data <= 11'd0;
end
//----------------------------��������----------------------
always @(*) begin
    if(!rst_n)
        image_data = 8'h0;
    else begin
        case(curr_state)
            HEAD_PACKET:begin
                case(cnt_data)                             
                    4'd0:image_data = HEAD[31:24];           
                    4'd1:image_data = HEAD[23:16];  
					4'd2:image_data = HEAD[15:8] ;           
                    4'd3:image_data = HEAD[7:0]  ;
					4'd4:image_data = ADDR;	
                    4'd5:image_data = DATA_NUM[31:24];
                    4'd6:image_data = DATA_NUM[23:16];
					4'd7:image_data = DATA_NUM[15:8];       
                    4'd8:image_data = DATA_NUM[7:0];  
					4'd9:image_data = CMD;   
                    default:image_data = cam_data; 
                endcase
            end
            DATA_PACKET:image_data = cam_data;
            LAST_PACKET:begin
                if(cnt_data == h_num)
                    image_data = CRC[15:8];
				else if(cnt_data == h_num + 16'd1)
					image_data = CRC[7:0];
                else 
                    image_data = cam_data;
            end
            default:image_data = 8'h0;
        endcase
    end
end
//----------------------------ddr��fifoʹ��----------------------
// always @(posedge clk or negedge rst_n) begin
    // if(!rst_n)
        // rf_rd_en <= 1'b0;
    // else if(udp_data_valid && ((curr_state == HEAD_PACKET && cnt_data >= 11'd9) || curr_state == DATA_PACKET || (curr_state == LAST_PACKET && cnt_data < h_num - 1)))
        // rf_rd_en <= 1'b1;
    // else
        // rf_rd_en <= 1'b0;
// end
assign rf_rd_en = udp_data_valid && 
                  ( (curr_state == HEAD_PACKET && cnt_data > 11'd8 && cnt_data < 11'd1289) || 
                    (curr_state == DATA_PACKET && cnt_data < h_num - 11'd1) || 
                    (curr_state == LAST_PACKET && cnt_data < h_num - 11'd1) 
                  );
//----------------------------��̫����ʼ�����ź�----------------------
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        udp_tx_data_start <= 1'b0;
    else if((next_state == HEAD_PACKET || next_state == DATA_PACKET || next_state == LAST_PACKET) && (curr_state != next_state))
        udp_tx_data_start <= 1'b1;
    else
        udp_tx_data_start <= 1'b0;
end
//----------------------------һ֡ͼ���͵ĸ���----------------------
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        cnt_h <= 11'd0;
    else if(curr_state == IDLE)
        cnt_h <= 11'd0;
    else if(udp_tx_done)
        cnt_h <= cnt_h + 11'd1;
    else
        cnt_h <= cnt_h;
end
//----------------------------��̫�������������ݸ���----------------------
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        image_data_num <= 16'd0;
    else if(curr_state == HEAD_PACKET)
        image_data_num <= h_num + 16'd10;
    else if(curr_state == DATA_PACKET)
        image_data_num <= h_num;
    else if(curr_state == LAST_PACKET)
        image_data_num <= h_num + 16'd2;
    else
        image_data_num <= image_data_num;
end

endmodule
