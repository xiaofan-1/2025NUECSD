module number_rom( 
	input	wire			clk				,
	input	wire			rst_n			,
	input	wire 	[11:0]  pixel_x			,
	input	wire 	[11:0]	pixel_y			,
	input	wire			de				,
	input	wire	[ 3:0]	number_data		,
    output 	reg  	[23:0] 	data_o		
);

reg  [511:0] char_num [9:0] ;  

reg 	[11:0]	addra;
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        addra <= 0;
    else if(addra == 512 - 1)
        addra <= 0;
    else if(addra < 512  && pixel_x < 16  && pixel_y < 82 && pixel_y > 50 && de)
        addra <= addra + 1;
end

always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        data_o <= 0;
    else if(char_num[number_data][addra] == 0)
        data_o <= 24'hff_ff_ff;
	else
		data_o <= 24'h0;
end

always @(posedge clk) begin 
    char_num[0] <= 512'h00000000000000000000000003C006200C30181818181808300C300C300C300C300C300C300C300C300C300C1808181818180C30062003C00000000000000000;/*"0",0*/
    char_num[1] <= 512'h000000000000000000000000008001801F800180018001800180018001800180018001800180018001800180018001800180018003C01FF80000000000000000;/*"1",1*/
    char_num[2] <= 512'h00000000000000000000000007E008381018200C200C300C300C000C001800180030006000C0018003000200040408041004200C3FF83FF80000000000000000;/*"2",2*/
    char_num[3] <= 512'h00000000000000000000000007C018603030301830183018001800180030006003C0007000180008000C000C300C300C30083018183007C00000000000000000;/*"3",3*/
    char_num[4] <= 512'h0000000000000000000000000060006000E000E0016001600260046004600860086010603060206040607FFC0060006000600060006003FC0000000000000000;/*"4",4*/
    char_num[5] <= 512'h0000000000000000000000000FFC0FFC10001000100010001000100013E0143018181008000C000C000C000C300C300C20182018183007C00000000000000000;/*"5",5*/
    char_num[6] <= 512'h00000000000000000000000001E006180C180818180010001000300033E0363038183808300C300C300C300C300C180C18080C180E3003E00000000000000000;/*"6",6*/
    char_num[7] <= 512'h0000000000000000000000001FFC1FFC100830102010202000200040004000400080008001000100010001000300030003000300030003000000000000000000;/*"7",7*/
    char_num[8] <= 512'h00000000000000000000000007E00C301818300C300C300C380C38081E180F2007C018F030783038601C600C600C600C600C3018183007C00000000000000000;/*"8",8*/
    char_num[9] <= 512'h00000000000000000000000007C01820301030186008600C600C600C600C600C701C302C186C0F8C000C0018001800103030306030C00F800000000000000000;/*"9",9*/
end

endmodule
